`timescale 10ns/1ns
`include "while_ex.v"

module while_ex_tb;
    /* // instantiate the module under test
    Repeat uut();
    $dumpfile("while_ex.vcd"); 
   // while_ex uut(); */


endmodule
